package router_pkg;

  import uvm_pkg::*;

  `include "uvm_macros.svh"

  `include "source_xtn.sv"
  `include "dest_xtn.sv"

  `include "source_config.sv"
  `include "dest_config.sv"
  `include "env_config.sv"

  `include "source_seqs.sv"
  `include "dest_seqs.sv"

  `include "source_drv.sv"
  `include "source_mon.sv"
  `include "source_sequencer.sv"
  `include "source_agent.sv"
  `include "source_agent_top.sv"

  `include "dest_drv.sv"
  `include "dest_mon.sv"
  `include "dest_sequencer.sv"
  `include "dest_agent.sv"
  `include "dest_agent_top.sv"

  `include "virtual_sequencer.sv"
  `include "virtual_seqs.sv"
  `include "scoreboard.sv"

  `include "env.sv"

  `include "base_test.sv"

endpackage


